library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity instructionMemory is
    port(
        clk : in std_logic;
        address : in std_logic_vector(15 downto 0);
        instruction : out std_logic_vector(15 downto 0)
    );
end entity instructionMemory;

architecture instructions of instructionMemory is
    type instructionMemoryDataType is array (0 to 127) of std_logic_vector(15 downto 0);
    signal instructionMemoryData : instructionMemoryDataType := (
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111", 
"1111111111111111"      
    );
begin 
    process(clk)
        begin
            if clk = '1' and clk'event then
                instruction <= instructionMemoryData(to_integer(unsigned(address)));
            end if;
    end process;
end architecture instructions;